entity top 