entity top a