LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE work.aux_package.all;
-------------------------------------------------------------
entity Datapath is
	generic (n : positive := 8 );
	port(
		clk : in std_logic;
		OPCin,OPC2,OPC1,Ld,Bin,Cout : in std_logic;
		DATAin  : in std_logic_vector(n-1 downto 0);
		---------------------------------------------
		Input,One : out std_logic;
		DATAout : out std_logic_vector(n-1 downto 0)
	);
end Datapath;
------------- complete the Datapath Unit Architecture code --------------
architecture arc_sys of Datapath is
signal reg_c,reg_b,ALUout,counter,one_before_not:STD_LOGIC_VECTOR(n-1 downto 0);
signal addersub_result,logical_result:STD_LOGIC_VECTOR(n-1 downto 0);
signal reg_opc,ALUFN:STD_LOGIC_VECTOR(2 downto 0); 
signal enable_dec,A,ctr_input std_logic;
alias Opcode :std_logic_vector(2 downto 0) is DATAin(2 downto 0);
);
begin
	ctr_input<= and DATAin ;
	ALUFN<= reg_opc when(OPC2='1') else "ZZZ";
	A<='1' when (OPC1='1') else 'Z';
	one_before_not(0) <= not counter(0);
	create_one:	for i in 1 to n-1 generate
		one_before_not(i) <= counter(i);
end generate;
	One <= nor one_before_not);

------------------------counter process--------------------------
d_counter : process(clk)
begin
	if (clk'event and clk='1') then -- rising edge
		if (Ld ='1') then
			counter <=DATAin;
		elsif (Ld ='0') then
			counter <= counter -1;
		end if;	
	end if;
end process;
------------------------Registers process--------------------------
reg_opc_proc : process(clk)
begin
	if (clk'event and clk='1') then -- rising edge
		if (OPCin='1') --register OPC
			reg_opc <= Opcode;
		end if;
		if (Bin='1') --register B
			reg_b <= ALUout;
		end if;
		if (Cout='1') --register C
			DATAout < =reg_c; -- out
		else
			reg_c<= reg_b; --in every operation cycle
		end if;
	end if;
end process;
-----------------------AdderSub---------------------------
AdderSubaba : AdderSub generic map (n)port map(
			sctr => ALUFN(1), --'1' SUB , '0' ADD
			x => DATAin,
			y => reg_b,
			s => addersub_result);	
-----------------------Logical----------------------------			
Logiloko : Logical generic map (n) port map( -- x and y are crossed twice duo to a loko programmer
			ALUFN => ALUFN(1 downto 0),
			x => DATAin,
			y => reg_b,
			result => logical_result);
-----------------------ALU--------------------------------					
ALUFORU  : ALU generic map (n) port map(
			ALUFN => ALUFN(2 downto 0), 
			--ALUFN := [0,0,0]=A ,[0,0,1]=A+B, [0,1,0]=A-B, [0,1,1]=AorB, [1,0,0]= AandB, [1,0,1]=AxorB 
			A => A,
			vector_A => DATAin,
			logical => logical_result
			addersub => addersub_result,
			ALUout=>ALUout);
end arc_sys;







